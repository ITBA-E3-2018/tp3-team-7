module ej1a(clk, I, S, B1, B2);
	

endmodule
